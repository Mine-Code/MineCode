module types

pub struct Program {
	do_once bool
}
